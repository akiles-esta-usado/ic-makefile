** sch_path: /workspaces/ic-makefile/samples/pmos1f/symbol/pmos1f.sch
.subckt pmos1f S G D B
*.PININFO S:B G:B D:B B:B
M1 D G S B pfet_03v3 L=0.28u W=0.42u nf=1 m=1
.ends
.end
