** sch_path: /workspaces/ic-makefile/samples/inv_sample/test/inv_sample_test.sch

.include /home/designer/.volare/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /home/designer/.volare/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical
.lib /home/designer/.volare/gf180mcuD/libs.tech/ngspice/sm141064.ngspice mimcap_statistical
.lib /home/designer/.volare/gf180mcuD/libs.tech/ngspice/sm141064.ngspice cap_mim
.lib /home/designer/.volare/gf180mcuD/libs.tech/ngspice/sm141064.ngspice res_typical
.lib /home/designer/.volare/gf180mcuD/libs.tech/ngspice/sm141064.ngspice bjt_typical
.lib /home/designer/.volare/gf180mcuD/libs.tech/ngspice/sm141064.ngspice moscap_typical


.control
write
set appendwrite
.endc


**.subckt inv_sample_test
x1 vdd out in vss inv_sample
vvdd vdd GND 3.3
vin in GND pulse(0 3.3 100p 100p 1n 4n 10n)
vvss vss GND 0
**** begin user architecture code


.control
save in out out_pex time

tran 0.01n 100n
*plot in out out_pex

write
.endc




.control
save in out out_pex time

tran 0.01n 20n
*plot in out out_pex

write
.endc




*.include inv_sample_pex.spice
.include ../layout_pex/inv_sample_pex.spice
Xinv_pex  vdd out_pex in vss inv_sample_pex




.control
save in out out_pex

dc vin 0 3.3 0.001
*plot out vs in out_pex vs in

write
.endc


**** end user architecture code
**.ends

* expanding   symbol:  symbol/inv_sample.sym # of pins=4
** sym_path: /workspaces/ic-makefile/samples/inv_sample/symbol/inv_sample.sym
** sch_path: /workspaces/ic-makefile/samples/inv_sample/symbol/inv_sample.sch
.subckt inv_sample vdd out in vss
*.iopin vdd
*.iopin out
*.iopin vss
*.iopin in
XM1 out in vdd vdd pfet_03v3 L=0.28u W=1.26u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
XM2 out in vss vss nfet_03v3 L=0.28u W=0.42u nf=1 ad='int((nf+1)/2) * W/nf * 0.18u' as='int((nf+2)/2) * W/nf * 0.18u' pd='2*int((nf+1)/2) * (W/nf + 0.18u)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.18u)' nrd='0.18u / W' nrs='0.18u / W' sa=0 sb=0 sd=0 m=1
.ends

.GLOBAL GND
.end
