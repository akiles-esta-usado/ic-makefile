* NGSPICE file created from sigma_delta_counter.ext - technology: sky130A

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_2 abstract view
.subckt sky130_fd_sc_hd__dfxtp_2 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

.subckt sigma_delta_counter VGND VPWR clk ones[0] ones[1] ones[2] ones[3] ones[4]
+ ones[5] ones[6] ones[7] ones[8] ones[9] pulse ready rst
XFILLER_0_13_73 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_131_ _074_ _069_ _075_ VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__and3b_1
XFILLER_0_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_114_ _060_ _062_ _058_ _063_ _039_ VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__o311a_1
Xoutput7 net7 VGND VGND VPWR VPWR ones[4] sky130_fd_sc_hd__buf_1
XFILLER_0_7_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_130_ net6 net5 _067_ net7 VGND VGND VPWR VPWR _075_ sky130_fd_sc_hd__a31o_1
XTAP_TAPCELL_ROW_8_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_113_ counter\[7\] counter\[8\] _054_ counter\[9\] VGND VGND VPWR VPWR _063_ sky130_fd_sc_hd__a31o_1
Xoutput10 net10 VGND VGND VPWR VPWR ones[7] sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput8 net8 VGND VGND VPWR VPWR ones[5] sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_2_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_8_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_112_ counter\[9\] VGND VGND VPWR VPWR _062_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_15_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput9 net9 VGND VGND VPWR VPWR ones[6] sky130_fd_sc_hd__buf_1
Xoutput11 net11 VGND VGND VPWR VPWR ones[8] sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_2_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_12_Left_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_111_ _060_ _058_ _061_ VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput12 net12 VGND VGND VPWR VPWR ones[9] sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_15_Left_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_0_Left_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_110_ counter\[7\] counter\[8\] _054_ _038_ net2 VGND VGND VPWR VPWR _061_ sky130_fd_sc_hd__a311o_1
XTAP_TAPCELL_ROW_15_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput13 net13 VGND VGND VPWR VPWR ready sky130_fd_sc_hd__buf_1
XFILLER_0_13_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_169_ clknet_1_1__leaf_clk _017_ VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__dfxtp_1
XFILLER_0_7_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_099_ _051_ _039_ _052_ VGND VGND VPWR VPWR _053_ sky130_fd_sc_hd__and3b_1
X_168_ clknet_1_0__leaf_clk _016_ VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_167_ clknet_1_1__leaf_clk _015_ VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__dfxtp_1
X_098_ counter\[4\] _047_ counter\[5\] VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__a21o_1
XPHY_EDGE_ROW_7_Left_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_7_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_166_ clknet_1_1__leaf_clk _014_ VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__dfxtp_1
X_097_ counter\[4\] counter\[5\] _047_ VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__and3_1
X_149_ _032_ _029_ _033_ VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_148_ net12 net11 _028_ net2 net13 VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__a311o_1
X_096_ _050_ VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__clkbuf_1
X_165_ clknet_1_0__leaf_clk _013_ VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__dfxtp_2
XTAP_TAPCELL_ROW_6_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_079_ counter\[3\] _035_ _036_ _037_ VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__and4b_1
XFILLER_0_7_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_164_ clknet_1_1__leaf_clk _012_ VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__dfxtp_1
X_095_ _048_ _039_ _049_ VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__and3b_1
XFILLER_0_10_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_078_ counter\[4\] counter\[5\] counter\[8\] counter\[9\] VGND VGND VPWR VPWR _037_
+ sky130_fd_sc_hd__and4b_1
X_147_ net12 VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_094_ counter\[4\] _047_ VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__nand2_1
X_163_ clknet_1_0__leaf_clk _011_ VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__dfxtp_1
X_077_ counter\[7\] counter\[6\] VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_11_Left_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_129_ net7 net6 _071_ VGND VGND VPWR VPWR _074_ sky130_fd_sc_hd__and3_1
X_146_ _031_ VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__buf_1
XFILLER_0_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_14_Left_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_162_ clknet_1_0__leaf_clk _010_ VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__dfxtp_2
X_093_ counter\[4\] _047_ VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_076_ counter\[0\] counter\[1\] counter\[2\] VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__and3_1
X_145_ _069_ _029_ _030_ VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__and3_1
Xinput1 pulse VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_128_ net6 _071_ _073_ VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_161_ clknet_1_1__leaf_clk _009_ VGND VGND VPWR VPWR counter\[9\] sky130_fd_sc_hd__dfxtp_1
X_092_ counter\[0\] counter\[1\] counter\[3\] counter\[2\] VGND VGND VPWR VPWR _047_
+ sky130_fd_sc_hd__and4_2
Xinput2 rst VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_2
X_127_ net6 _071_ _069_ VGND VGND VPWR VPWR _073_ sky130_fd_sc_hd__o21ai_1
X_144_ _024_ _027_ net11 VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_143_ net11 _028_ VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__nand2_1
XFILLER_0_11_76 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_160_ clknet_1_0__leaf_clk _008_ VGND VGND VPWR VPWR counter\[8\] sky130_fd_sc_hd__dfxtp_1
X_091_ _046_ VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__clkbuf_1
X_126_ net5 _067_ _069_ _072_ VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_109_ counter\[8\] VGND VGND VPWR VPWR _060_ sky130_fd_sc_hd__inv_2
X_090_ _039_ _045_ VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_9_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_3_Left_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_125_ _071_ VGND VGND VPWR VPWR _072_ sky130_fd_sc_hd__inv_2
X_142_ _026_ _025_ _028_ net13 net2 VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__a2111oi_1
XPHY_EDGE_ROW_6_Left_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_108_ _059_ VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_3_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_141_ net6 _071_ _023_ _027_ VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_10_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_124_ net5 net4 net3 net1 VGND VGND VPWR VPWR _071_ sky130_fd_sc_hd__and4_2
X_107_ _039_ _057_ _058_ VGND VGND VPWR VPWR _059_ sky130_fd_sc_hd__and3_1
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_140_ net10 net9 VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__and2_1
X_106_ counter\[7\] _054_ VGND VGND VPWR VPWR _058_ sky130_fd_sc_hd__nand2_1
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_123_ _067_ _070_ VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_122_ net4 _068_ _069_ VGND VGND VPWR VPWR _070_ sky130_fd_sc_hd__o21ai_1
XTAP_TAPCELL_ROW_4_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_105_ counter\[7\] _054_ VGND VGND VPWR VPWR _057_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_12 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_11_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_121_ net13 net2 VGND VGND VPWR VPWR _069_ sky130_fd_sc_hd__nor2_2
XPHY_EDGE_ROW_10_Left_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_104_ _056_ VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_1_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_14_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_24 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_120_ net13 net1 net3 VGND VGND VPWR VPWR _068_ sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_49 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_103_ _054_ _039_ _055_ VGND VGND VPWR VPWR _056_ sky130_fd_sc_hd__and3b_1
XFILLER_0_8_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_102_ counter\[6\] _051_ VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_101_ counter\[4\] counter\[5\] counter\[6\] _047_ VGND VGND VPWR VPWR _054_ sky130_fd_sc_hd__and4_2
XFILLER_0_3_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_2_Left_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_100_ _053_ VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_7_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_5_Left_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_159_ clknet_1_1__leaf_clk _007_ VGND VGND VPWR VPWR counter\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_158_ clknet_1_1__leaf_clk _006_ VGND VGND VPWR VPWR counter\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_089_ counter\[3\] _035_ VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__xor2_1
XFILLER_0_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_1_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_1_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_9_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_088_ net2 _035_ _044_ VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__nor3_1
X_157_ clknet_1_0__leaf_clk _005_ VGND VGND VPWR VPWR counter\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_9_Left_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_156_ clknet_1_1__leaf_clk _004_ VGND VGND VPWR VPWR counter\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_087_ counter\[0\] counter\[1\] counter\[2\] VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__a21oi_1
X_139_ net10 VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_6 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_086_ _043_ VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__clkbuf_1
X_155_ clknet_1_0__leaf_clk _003_ VGND VGND VPWR VPWR counter\[3\] sky130_fd_sc_hd__dfxtp_1
X_172_ clknet_1_0__leaf_clk _020_ VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__dfxtp_2
X_138_ net9 _024_ _025_ _069_ VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__o211a_1
XFILLER_0_0_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_4_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_171_ clknet_1_0__leaf_clk _019_ VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__dfxtp_1
X_154_ clknet_1_1__leaf_clk _002_ VGND VGND VPWR VPWR counter\[2\] sky130_fd_sc_hd__dfxtp_1
X_085_ _041_ _039_ _042_ VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__and3_1
XFILLER_0_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_137_ net9 net8 _074_ VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__nand3_1
XFILLER_0_9_10 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_170_ clknet_1_1__leaf_clk _018_ VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_13_Left_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_084_ counter\[0\] counter\[1\] VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__or2_1
X_136_ net6 net5 _067_ _023_ VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__and4_1
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_153_ clknet_1_0__leaf_clk _001_ VGND VGND VPWR VPWR counter\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_15_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_119_ net13 net1 net4 net3 VGND VGND VPWR VPWR _067_ sky130_fd_sc_hd__o211a_1
XPHY_EDGE_ROW_1_Left_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_152_ clknet_1_1__leaf_clk _000_ VGND VGND VPWR VPWR counter\[0\] sky130_fd_sc_hd__dfxtp_1
X_083_ counter\[0\] counter\[1\] VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__nand2_1
XFILLER_0_3_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_135_ net8 net7 VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_78 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_4_Left_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_118_ _065_ _066_ VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput3 net3 VGND VGND VPWR VPWR ones[0] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_151_ _034_ VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_134_ net8 _074_ _022_ VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__a21oi_1
X_082_ _040_ VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_117_ net3 _064_ net1 net2 VGND VGND VPWR VPWR _066_ sky130_fd_sc_hd__a31o_1
XFILLER_0_12_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput4 net4 VGND VGND VPWR VPWR ones[1] sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_12_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_081_ counter\[0\] _039_ VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__and2b_1
X_150_ net2 _038_ VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__and2b_1
XFILLER_0_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_133_ net8 _074_ _069_ VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_116_ net3 _064_ net1 VGND VGND VPWR VPWR _065_ sky130_fd_sc_hd__a21oi_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput5 net5 VGND VGND VPWR VPWR ones[2] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_080_ net2 _038_ VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__nor2_2
X_132_ _021_ VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Left_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_115_ net13 VGND VGND VPWR VPWR _064_ sky130_fd_sc_hd__inv_2
Xoutput6 net6 VGND VGND VPWR VPWR ones[3] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
.ends

